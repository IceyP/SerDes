library verilog;
use verilog.vl_types.all;
entity tg is
    generic(
        C_AXI_ADDR_WIDTH: integer := 32;
        C_AXI_DATA_WIDTH: integer := 32;
        C_AXI_NBURST_SUPPORT: integer := 0;
        C_BEGIN_ADDRESS : integer := 0;
        C_END_ADDRESS   : integer := 255;
        C_EN_WRAP_TRANS : integer := 0;
        CTL_SIG_WIDTH   : integer := 3;
        WR_STS_WIDTH    : integer := 16;
        RD_STS_WIDTH    : integer := 16;
        DBG_WR_STS_WIDTH: integer := 32;
        DBG_RD_STS_WIDTH: integer := 32;
        ENFORCE_RD_WR   : integer := 0;
        ENFORCE_RD_WR_CMD: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        ENFORCE_RD_WR_PATTERN: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0)
    );
    port(
        clk             : in     vl_logic;
        resetn          : in     vl_logic;
        init_cmptd      : in     vl_logic;
        init_test       : in     vl_logic;
        wrap_en         : in     vl_logic;
        cmd_ack         : in     vl_logic;
        cmd_en          : out    vl_logic;
        cmd             : out    vl_logic_vector(2 downto 0);
        blen            : out    vl_logic_vector(7 downto 0);
        addr            : out    vl_logic_vector(31 downto 0);
        ctl             : out    vl_logic_vector;
        wdata_rdy       : in     vl_logic;
        wdata_vld       : out    vl_logic;
        wdata_cmptd     : out    vl_logic;
        wdata           : out    vl_logic_vector;
        wdata_bvld      : out    vl_logic_vector;
        wdata_sts_vld   : in     vl_logic;
        wdata_sts       : in     vl_logic_vector;
        rdata_vld       : in     vl_logic;
        rdata           : in     vl_logic_vector;
        rdata_bvld      : in     vl_logic_vector;
        rdata_cmptd     : in     vl_logic;
        rdata_sts       : in     vl_logic_vector;
        rdata_rdy       : out    vl_logic;
        cmd_err         : out    vl_logic;
        data_msmatch_err: out    vl_logic;
        write_err       : out    vl_logic;
        read_err        : out    vl_logic;
        test_cmptd      : out    vl_logic;
        write_cmptd     : out    vl_logic;
        read_cmptd      : out    vl_logic;
        cmptd_cycle     : out    vl_logic;
        dbg_wr_sts_vld  : out    vl_logic;
        dbg_wr_sts      : out    vl_logic_vector;
        dbg_rd_sts_vld  : out    vl_logic;
        dbg_rd_sts      : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of C_AXI_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_AXI_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_AXI_NBURST_SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of C_BEGIN_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of C_END_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of C_EN_WRAP_TRANS : constant is 1;
    attribute mti_svvh_generic_type of CTL_SIG_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of WR_STS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of RD_STS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DBG_WR_STS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DBG_RD_STS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ENFORCE_RD_WR : constant is 1;
    attribute mti_svvh_generic_type of ENFORCE_RD_WR_CMD : constant is 1;
    attribute mti_svvh_generic_type of ENFORCE_RD_WR_PATTERN : constant is 1;
end tg;
