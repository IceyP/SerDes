---------------------------------------------------------------------
--                   Auto gen By QAMmap                            --
--  For QAM 256 input format is 1xxxxxx                            --
--  For QAM 128 input format is 01xxxxx                            --
--  For QAM  64 input format is 001xxxx                            --
--  For QAM  32 input format is 0001xxx                            --
--  For QAM  16 input format is 00001xx                            --
--  Output is I/Q 4bit without sign                                --
---------------------------------------------------------------------
library IEEE;                                                        
use IEEE.STD_LOGIC_1164.all;                                         
                                                                     
entity QAMRom is                                                     
	 port(  
         clk : in STD_LOGIC;
		 rst : in std_logic; 
		 D : in STD_LOGIC_VECTOR(6 downto 0);                            
		 I : out STD_LOGIC_VECTOR(3 downto 0);                           
		 Q : out STD_LOGIC_VECTOR(3 downto 0)                            
	     );                                                            
end QAMRom;                                                          
                                                                     
architecture behave of QAMRom is                                     
                                                                     
begin                                                                
                                                                     
IRom : process(clk,rst)                                                 
begin 
    if rst='1' then
        I <= "0000";
	elsif rising_edge(clk) then
        case D is                                                        
        when "0000100" => I<="0001";
        when "0000101" => I<="0011";
        when "0000110" => I<="0001";
        when "0000111" => I<="0011";
        when "0001000" => I<="0001";
        when "0001001" => I<="0011";
        when "0001011" => I<="0101";
        when "0001100" => I<="0001";
        when "0001101" => I<="0011";
        when "0001111" => I<="0101";
        when "0001110" => I<="0001";
        when "0001010" => I<="0011";
        when "0010000" => I<="0001";
        when "0010001" => I<="0011";
        when "0010101" => I<="0101";
        when "0010100" => I<="0111";
        when "0010010" => I<="0001";
        when "0010011" => I<="0011";
        when "0010111" => I<="0101";
        when "0010110" => I<="0111";
        when "0011010" => I<="0001";
        when "0011011" => I<="0011";
        when "0011111" => I<="0101";
        when "0011110" => I<="0111";
        when "0011000" => I<="0001";
        when "0011001" => I<="0011";
        when "0011101" => I<="0101";
        when "0011100" => I<="0111";
        when "0100000" => I<="0001";
        when "0100001" => I<="0011";
        when "0100101" => I<="0101";
        when "0100100" => I<="0111";
        when "0101100" => I<="1001";
        when "0101101" => I<="1011";
        when "0100010" => I<="0001";
        when "0100011" => I<="0011";
        when "0100111" => I<="0101";
        when "0100110" => I<="0111";
        when "0101110" => I<="1001";
        when "0101111" => I<="1011";
        when "0110010" => I<="0001";
        when "0110011" => I<="0011";
        when "0110111" => I<="0101";
        when "0110110" => I<="0111";
        when "0111110" => I<="1001";
        when "0111111" => I<="1011";
        when "0110000" => I<="0001";
        when "0110001" => I<="0011";
        when "0110101" => I<="0101";
        when "0110100" => I<="0111";
        when "0111100" => I<="1001";
        when "0111101" => I<="1011";
        when "0111000" => I<="0001";
        when "0111001" => I<="0011";
        when "0101001" => I<="0101";
        when "0101000" => I<="0111";
        when "0111010" => I<="0001";
        when "0111011" => I<="0011";
        when "0101011" => I<="0101";
        when "0101010" => I<="0111";
        when "1000000" => I<="0001";
        when "1000001" => I<="0011";
        when "1000101" => I<="0101";
        when "1000100" => I<="0111";
        when "1010100" => I<="1001";
        when "1010101" => I<="1011";
        when "1010001" => I<="1101";
        when "1010000" => I<="1111";
        when "1000010" => I<="0001";
        when "1000011" => I<="0011";
        when "1000111" => I<="0101";
        when "1000110" => I<="0111";
        when "1010110" => I<="1001";
        when "1010111" => I<="1011";
        when "1010011" => I<="1101";
        when "1010010" => I<="1111";
        when "1001010" => I<="0001";
        when "1001011" => I<="0011";
        when "1001111" => I<="0101";
        when "1001110" => I<="0111";
        when "1011110" => I<="1001";
        when "1011111" => I<="1011";
        when "1011011" => I<="1101";
        when "1011010" => I<="1111";
        when "1001000" => I<="0001";
        when "1001001" => I<="0011";
        when "1001101" => I<="0101";
        when "1001100" => I<="0111";
        when "1011100" => I<="1001";
        when "1011101" => I<="1011";
        when "1011001" => I<="1101";
        when "1011000" => I<="1111";
        when "1101000" => I<="0001";
        when "1101001" => I<="0011";
        when "1101101" => I<="0101";
        when "1101100" => I<="0111";
        when "1111100" => I<="1001";
        when "1111101" => I<="1011";
        when "1111001" => I<="1101";
        when "1111000" => I<="1111";
        when "1101010" => I<="0001";
        when "1101011" => I<="0011";
        when "1101111" => I<="0101";
        when "1101110" => I<="0111";
        when "1111110" => I<="1001";
        when "1111111" => I<="1011";
        when "1111011" => I<="1101";
        when "1111010" => I<="1111";
        when "1100010" => I<="0001";
        when "1100011" => I<="0011";
        when "1100111" => I<="0101";
        when "1100110" => I<="0111";
        when "1110110" => I<="1001";
        when "1110111" => I<="1011";
        when "1110011" => I<="1101";
        when "1110010" => I<="1111";
        when "1100000" => I<="0001";
        when "1100001" => I<="0011";
        when "1100101" => I<="0101";
        when "1100100" => I<="0111";
        when "1110100" => I<="1001";
        when "1110101" => I<="1011";
        when "1110001" => I<="1101";
        when "1110000" => I<="1111";
        when others => I<=( others=>'0' );                           
        end case;
    end if;	
end process;                                                         
                                                                     
QRom : process(clk,rst)                                                 
begin 
    if rst='1' then
        Q <= "0000";
	elsif rising_edge(clk) then                                                                
        case D is                                                       
        when "0000100" => Q<="0001";
        when "0000101" => Q<="0001";
        when "0000110" => Q<="0011";
        when "0000111" => Q<="0011";
        when "0001000" => Q<="0001";
        when "0001001" => Q<="0001";
        when "0001011" => Q<="0001";
        when "0001100" => Q<="0011";
        when "0001101" => Q<="0011";
        when "0001111" => Q<="0011";
        when "0001110" => Q<="0101";
        when "0001010" => Q<="0101";
        when "0010000" => Q<="0001";
        when "0010001" => Q<="0001";
        when "0010101" => Q<="0001";
        when "0010100" => Q<="0001";
        when "0010010" => Q<="0011";
        when "0010011" => Q<="0011";
        when "0010111" => Q<="0011";
        when "0010110" => Q<="0011";
        when "0011010" => Q<="0101";
        when "0011011" => Q<="0101";
        when "0011111" => Q<="0101";
        when "0011110" => Q<="0101";
        when "0011000" => Q<="0111";
        when "0011001" => Q<="0111";
        when "0011101" => Q<="0111";
        when "0011100" => Q<="0111";
        when "0100000" => Q<="0001";
        when "0100001" => Q<="0001";
        when "0100101" => Q<="0001";
        when "0100100" => Q<="0001";
        when "0101100" => Q<="0001";
        when "0101101" => Q<="0001";
        when "0100010" => Q<="0011";
        when "0100011" => Q<="0011";
        when "0100111" => Q<="0011";
        when "0100110" => Q<="0011";
        when "0101110" => Q<="0011";
        when "0101111" => Q<="0011";
        when "0110010" => Q<="0101";
        when "0110011" => Q<="0101";
        when "0110111" => Q<="0101";
        when "0110110" => Q<="0101";
        when "0111110" => Q<="0101";
        when "0111111" => Q<="0101";
        when "0110000" => Q<="0111";
        when "0110001" => Q<="0111";
        when "0110101" => Q<="0111";
        when "0110100" => Q<="0111";
        when "0111100" => Q<="0111";
        when "0111101" => Q<="0111";
        when "0111000" => Q<="1001";
        when "0111001" => Q<="1001";
        when "0101001" => Q<="1001";
        when "0101000" => Q<="1001";
        when "0111010" => Q<="1011";
        when "0111011" => Q<="1011";
        when "0101011" => Q<="1011";
        when "0101010" => Q<="1011";
        when "1000000" => Q<="0001";
        when "1000001" => Q<="0001";
        when "1000101" => Q<="0001";
        when "1000100" => Q<="0001";
        when "1010100" => Q<="0001";
        when "1010101" => Q<="0001";
        when "1010001" => Q<="0001";
        when "1010000" => Q<="0001";
        when "1000010" => Q<="0011";
        when "1000011" => Q<="0011";
        when "1000111" => Q<="0011";
        when "1000110" => Q<="0011";
        when "1010110" => Q<="0011";
        when "1010111" => Q<="0011";
        when "1010011" => Q<="0011";
        when "1010010" => Q<="0011";
        when "1001010" => Q<="0101";
        when "1001011" => Q<="0101";
        when "1001111" => Q<="0101";
        when "1001110" => Q<="0101";
        when "1011110" => Q<="0101";
        when "1011111" => Q<="0101";
        when "1011011" => Q<="0101";
        when "1011010" => Q<="0101";
        when "1001000" => Q<="0111";
        when "1001001" => Q<="0111";
        when "1001101" => Q<="0111";
        when "1001100" => Q<="0111";
        when "1011100" => Q<="0111";
        when "1011101" => Q<="0111";
        when "1011001" => Q<="0111";
        when "1011000" => Q<="0111";
        when "1101000" => Q<="1001";
        when "1101001" => Q<="1001";
        when "1101101" => Q<="1001";
        when "1101100" => Q<="1001";
        when "1111100" => Q<="1001";
        when "1111101" => Q<="1001";
        when "1111001" => Q<="1001";
        when "1111000" => Q<="1001";
        when "1101010" => Q<="1011";
        when "1101011" => Q<="1011";
        when "1101111" => Q<="1011";
        when "1101110" => Q<="1011";
        when "1111110" => Q<="1011";
        when "1111111" => Q<="1011";
        when "1111011" => Q<="1011";
        when "1111010" => Q<="1011";
        when "1100010" => Q<="1101";
        when "1100011" => Q<="1101";
        when "1100111" => Q<="1101";
        when "1100110" => Q<="1101";
        when "1110110" => Q<="1101";
        when "1110111" => Q<="1101";
        when "1110011" => Q<="1101";
        when "1110010" => Q<="1101";
        when "1100000" => Q<="1111";
        when "1100001" => Q<="1111";
        when "1100101" => Q<="1111";
        when "1100100" => Q<="1111";
        when "1110100" => Q<="1111";
        when "1110101" => Q<="1111";
        when "1110001" => Q<="1111";
        when "1110000" => Q<="1111";
        when others => Q<=( others=>'0' );                           
        end case; 
    end if;		
end process;                                                         
                                                                     
end behave;                                                          
