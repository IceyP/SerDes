library verilog;
use verilog.vl_types.all;
entity s6_axi4_tg is
    generic(
        C_PORT_CONFIG   : string  := "B32_B32_W32_R32_W32_R32";
        C_P0_PORT_MODE  : string  := "BI_MODE";
        C_P1_PORT_MODE  : string  := "BI_MODE";
        C_P2_PORT_MODE  : string  := "WR_MODE";
        C_P3_PORT_MODE  : string  := "RD_MODE";
        C_P4_PORT_MODE  : string  := "WR_MODE";
        C_P5_PORT_MODE  : string  := "RD_MODE";
        C_PORT_ENABLE   : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        C_BEGIN_ADDRESS : integer := 256;
        C_END_ADDRESS   : integer := 767;
        C_PRBS_EADDR_MASK_POS: vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        C_PRBS_SADDR_MASK_POS: integer := 256;
        C_EN_UPSIZER    : integer := 0;
        C_AXI_NBURST_SUPPORT: integer := 0;
        C_ENFORCE_RD_WR : integer := 0;
        C_ENFORCE_RD_WR_CMD: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        C_ENFORCE_RD_WR_PATTERN: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        C_EN_WRAP_TRANS : integer := 0;
        C_P0_AXI_SUPPORTS_READ: integer := 1;
        C_P0_AXI_SUPPORTS_WRITE: integer := 1;
        C_P0_AXI_ID_WIDTH: integer := 4;
        C_P0_AXI_ADDR_WIDTH: integer := 32;
        C_P0_AXI_DATA_WIDTH: integer := 32;
        C_P1_AXI_SUPPORTS_READ: integer := 1;
        C_P1_AXI_SUPPORTS_WRITE: integer := 1;
        C_P1_AXI_ID_WIDTH: integer := 4;
        C_P1_AXI_ADDR_WIDTH: integer := 32;
        C_P1_AXI_DATA_WIDTH: integer := 32;
        C_P2_AXI_SUPPORTS_READ: integer := 0;
        C_P2_AXI_SUPPORTS_WRITE: integer := 1;
        C_P2_AXI_ID_WIDTH: integer := 4;
        C_P2_AXI_ADDR_WIDTH: integer := 32;
        C_P2_AXI_DATA_WIDTH: integer := 32;
        C_P3_AXI_SUPPORTS_READ: integer := 1;
        C_P3_AXI_SUPPORTS_WRITE: integer := 0;
        C_P3_AXI_ID_WIDTH: integer := 4;
        C_P3_AXI_ADDR_WIDTH: integer := 32;
        C_P3_AXI_DATA_WIDTH: integer := 32;
        C_P4_AXI_SUPPORTS_READ: integer := 0;
        C_P4_AXI_SUPPORTS_WRITE: integer := 1;
        C_P4_AXI_ID_WIDTH: integer := 4;
        C_P4_AXI_ADDR_WIDTH: integer := 32;
        C_P4_AXI_DATA_WIDTH: integer := 32;
        C_P5_AXI_SUPPORTS_READ: integer := 1;
        C_P5_AXI_SUPPORTS_WRITE: integer := 0;
        C_P5_AXI_ID_WIDTH: integer := 4;
        C_P5_AXI_ADDR_WIDTH: integer := 32;
        C_P5_AXI_DATA_WIDTH: integer := 32;
        DBG_WR_STS_WIDTH: integer := 32;
        DBG_RD_STS_WIDTH: integer := 32
    );
    port(
        aclk            : in     vl_logic;
        aresetn         : in     vl_logic;
        init_cmptd      : in     vl_logic;
        init_test       : in     vl_logic;
        wdog_mask       : in     vl_logic;
        wrap_en         : in     vl_logic;
        axi_wready_c_p0 : in     vl_logic;
        axi_wid_c_p0    : out    vl_logic_vector;
        axi_waddr_c_p0  : out    vl_logic_vector;
        axi_wlen_c_p0   : out    vl_logic_vector(7 downto 0);
        axi_wsize_c_p0  : out    vl_logic_vector(2 downto 0);
        axi_wburst_c_p0 : out    vl_logic_vector(1 downto 0);
        axi_wlock_c_p0  : out    vl_logic;
        axi_wcache_c_p0 : out    vl_logic_vector(3 downto 0);
        axi_wprot_c_p0  : out    vl_logic_vector(2 downto 0);
        axi_wvalid_c_p0 : out    vl_logic;
        axi_wd_wready_c_p0: in     vl_logic;
        axi_wd_wid_c_p0 : out    vl_logic_vector;
        axi_wd_data_c_p0: out    vl_logic_vector;
        axi_wd_strb_c_p0: out    vl_logic_vector;
        axi_wd_last_c_p0: out    vl_logic;
        axi_wd_valid_c_p0: out    vl_logic;
        axi_wd_bid_c_p0 : in     vl_logic_vector;
        axi_wd_bresp_c_p0: in     vl_logic_vector(1 downto 0);
        axi_wd_bvalid_c_p0: in     vl_logic;
        axi_wd_bready_c_p0: out    vl_logic;
        axi_rready_c_p0 : in     vl_logic;
        axi_rid_c_p0    : out    vl_logic_vector;
        axi_raddr_c_p0  : out    vl_logic_vector;
        axi_rlen_c_p0   : out    vl_logic_vector(7 downto 0);
        axi_rsize_c_p0  : out    vl_logic_vector(2 downto 0);
        axi_rburst_c_p0 : out    vl_logic_vector(1 downto 0);
        axi_rlock_c_p0  : out    vl_logic;
        axi_rcache_c_p0 : out    vl_logic_vector(3 downto 0);
        axi_rprot_c_p0  : out    vl_logic_vector(2 downto 0);
        axi_rvalid_c_p0 : out    vl_logic;
        axi_rd_bid_c_p0 : in     vl_logic_vector;
        axi_rd_rresp_c_p0: in     vl_logic_vector(1 downto 0);
        axi_rd_rvalid_c_p0: in     vl_logic;
        axi_rd_data_c_p0: in     vl_logic_vector;
        axi_rd_last_c_p0: in     vl_logic;
        axi_rd_rready_c_p0: out    vl_logic;
        axi_wready_c_p1 : in     vl_logic;
        axi_wid_c_p1    : out    vl_logic_vector;
        axi_waddr_c_p1  : out    vl_logic_vector;
        axi_wlen_c_p1   : out    vl_logic_vector(7 downto 0);
        axi_wsize_c_p1  : out    vl_logic_vector(2 downto 0);
        axi_wburst_c_p1 : out    vl_logic_vector(1 downto 0);
        axi_wlock_c_p1  : out    vl_logic;
        axi_wcache_c_p1 : out    vl_logic_vector(3 downto 0);
        axi_wprot_c_p1  : out    vl_logic_vector(2 downto 0);
        axi_wvalid_c_p1 : out    vl_logic;
        axi_wd_wready_c_p1: in     vl_logic;
        axi_wd_wid_c_p1 : out    vl_logic_vector;
        axi_wd_data_c_p1: out    vl_logic_vector;
        axi_wd_strb_c_p1: out    vl_logic_vector;
        axi_wd_last_c_p1: out    vl_logic;
        axi_wd_valid_c_p1: out    vl_logic;
        axi_wd_bid_c_p1 : in     vl_logic_vector;
        axi_wd_bresp_c_p1: in     vl_logic_vector(1 downto 0);
        axi_wd_bvalid_c_p1: in     vl_logic;
        axi_wd_bready_c_p1: out    vl_logic;
        axi_rready_c_p1 : in     vl_logic;
        axi_rid_c_p1    : out    vl_logic_vector;
        axi_raddr_c_p1  : out    vl_logic_vector;
        axi_rlen_c_p1   : out    vl_logic_vector(7 downto 0);
        axi_rsize_c_p1  : out    vl_logic_vector(2 downto 0);
        axi_rburst_c_p1 : out    vl_logic_vector(1 downto 0);
        axi_rlock_c_p1  : out    vl_logic;
        axi_rcache_c_p1 : out    vl_logic_vector(3 downto 0);
        axi_rprot_c_p1  : out    vl_logic_vector(2 downto 0);
        axi_rvalid_c_p1 : out    vl_logic;
        axi_rd_bid_c_p1 : in     vl_logic_vector;
        axi_rd_rresp_c_p1: in     vl_logic_vector(1 downto 0);
        axi_rd_rvalid_c_p1: in     vl_logic;
        axi_rd_data_c_p1: in     vl_logic_vector;
        axi_rd_last_c_p1: in     vl_logic;
        axi_rd_rready_c_p1: out    vl_logic;
        axi_wready_c_p2 : in     vl_logic;
        axi_wid_c_p2    : out    vl_logic_vector;
        axi_waddr_c_p2  : out    vl_logic_vector;
        axi_wlen_c_p2   : out    vl_logic_vector(7 downto 0);
        axi_wsize_c_p2  : out    vl_logic_vector(2 downto 0);
        axi_wburst_c_p2 : out    vl_logic_vector(1 downto 0);
        axi_wlock_c_p2  : out    vl_logic;
        axi_wcache_c_p2 : out    vl_logic_vector(3 downto 0);
        axi_wprot_c_p2  : out    vl_logic_vector(2 downto 0);
        axi_wvalid_c_p2 : out    vl_logic;
        axi_wd_wready_c_p2: in     vl_logic;
        axi_wd_wid_c_p2 : out    vl_logic_vector;
        axi_wd_data_c_p2: out    vl_logic_vector;
        axi_wd_strb_c_p2: out    vl_logic_vector;
        axi_wd_last_c_p2: out    vl_logic;
        axi_wd_valid_c_p2: out    vl_logic;
        axi_wd_bid_c_p2 : in     vl_logic_vector;
        axi_wd_bresp_c_p2: in     vl_logic_vector(1 downto 0);
        axi_wd_bvalid_c_p2: in     vl_logic;
        axi_wd_bready_c_p2: out    vl_logic;
        axi_rready_c_p2 : in     vl_logic;
        axi_rid_c_p2    : out    vl_logic_vector;
        axi_raddr_c_p2  : out    vl_logic_vector;
        axi_rlen_c_p2   : out    vl_logic_vector(7 downto 0);
        axi_rsize_c_p2  : out    vl_logic_vector(2 downto 0);
        axi_rburst_c_p2 : out    vl_logic_vector(1 downto 0);
        axi_rlock_c_p2  : out    vl_logic;
        axi_rcache_c_p2 : out    vl_logic_vector(3 downto 0);
        axi_rprot_c_p2  : out    vl_logic_vector(2 downto 0);
        axi_rvalid_c_p2 : out    vl_logic;
        axi_rd_bid_c_p2 : in     vl_logic_vector;
        axi_rd_rresp_c_p2: in     vl_logic_vector(1 downto 0);
        axi_rd_rvalid_c_p2: in     vl_logic;
        axi_rd_data_c_p2: in     vl_logic_vector;
        axi_rd_last_c_p2: in     vl_logic;
        axi_rd_rready_c_p2: out    vl_logic;
        axi_wready_c_p3 : in     vl_logic;
        axi_wid_c_p3    : out    vl_logic_vector;
        axi_waddr_c_p3  : out    vl_logic_vector;
        axi_wlen_c_p3   : out    vl_logic_vector(7 downto 0);
        axi_wsize_c_p3  : out    vl_logic_vector(2 downto 0);
        axi_wburst_c_p3 : out    vl_logic_vector(1 downto 0);
        axi_wlock_c_p3  : out    vl_logic;
        axi_wcache_c_p3 : out    vl_logic_vector(3 downto 0);
        axi_wprot_c_p3  : out    vl_logic_vector(2 downto 0);
        axi_wvalid_c_p3 : out    vl_logic;
        axi_wd_wready_c_p3: in     vl_logic;
        axi_wd_wid_c_p3 : out    vl_logic_vector;
        axi_wd_data_c_p3: out    vl_logic_vector;
        axi_wd_strb_c_p3: out    vl_logic_vector;
        axi_wd_last_c_p3: out    vl_logic;
        axi_wd_valid_c_p3: out    vl_logic;
        axi_wd_bid_c_p3 : in     vl_logic_vector;
        axi_wd_bresp_c_p3: in     vl_logic_vector(1 downto 0);
        axi_wd_bvalid_c_p3: in     vl_logic;
        axi_wd_bready_c_p3: out    vl_logic;
        axi_rready_c_p3 : in     vl_logic;
        axi_rid_c_p3    : out    vl_logic_vector;
        axi_raddr_c_p3  : out    vl_logic_vector;
        axi_rlen_c_p3   : out    vl_logic_vector(7 downto 0);
        axi_rsize_c_p3  : out    vl_logic_vector(2 downto 0);
        axi_rburst_c_p3 : out    vl_logic_vector(1 downto 0);
        axi_rlock_c_p3  : out    vl_logic;
        axi_rcache_c_p3 : out    vl_logic_vector(3 downto 0);
        axi_rprot_c_p3  : out    vl_logic_vector(2 downto 0);
        axi_rvalid_c_p3 : out    vl_logic;
        axi_rd_bid_c_p3 : in     vl_logic_vector;
        axi_rd_rresp_c_p3: in     vl_logic_vector(1 downto 0);
        axi_rd_rvalid_c_p3: in     vl_logic;
        axi_rd_data_c_p3: in     vl_logic_vector;
        axi_rd_last_c_p3: in     vl_logic;
        axi_rd_rready_c_p3: out    vl_logic;
        axi_wready_c_p4 : in     vl_logic;
        axi_wid_c_p4    : out    vl_logic_vector;
        axi_waddr_c_p4  : out    vl_logic_vector;
        axi_wlen_c_p4   : out    vl_logic_vector(7 downto 0);
        axi_wsize_c_p4  : out    vl_logic_vector(2 downto 0);
        axi_wburst_c_p4 : out    vl_logic_vector(1 downto 0);
        axi_wlock_c_p4  : out    vl_logic;
        axi_wcache_c_p4 : out    vl_logic_vector(3 downto 0);
        axi_wprot_c_p4  : out    vl_logic_vector(2 downto 0);
        axi_wvalid_c_p4 : out    vl_logic;
        axi_wd_wready_c_p4: in     vl_logic;
        axi_wd_wid_c_p4 : out    vl_logic_vector;
        axi_wd_data_c_p4: out    vl_logic_vector;
        axi_wd_strb_c_p4: out    vl_logic_vector;
        axi_wd_last_c_p4: out    vl_logic;
        axi_wd_valid_c_p4: out    vl_logic;
        axi_wd_bid_c_p4 : in     vl_logic_vector;
        axi_wd_bresp_c_p4: in     vl_logic_vector(1 downto 0);
        axi_wd_bvalid_c_p4: in     vl_logic;
        axi_wd_bready_c_p4: out    vl_logic;
        axi_rready_c_p4 : in     vl_logic;
        axi_rid_c_p4    : out    vl_logic_vector;
        axi_raddr_c_p4  : out    vl_logic_vector;
        axi_rlen_c_p4   : out    vl_logic_vector(7 downto 0);
        axi_rsize_c_p4  : out    vl_logic_vector(2 downto 0);
        axi_rburst_c_p4 : out    vl_logic_vector(1 downto 0);
        axi_rlock_c_p4  : out    vl_logic;
        axi_rcache_c_p4 : out    vl_logic_vector(3 downto 0);
        axi_rprot_c_p4  : out    vl_logic_vector(2 downto 0);
        axi_rvalid_c_p4 : out    vl_logic;
        axi_rd_bid_c_p4 : in     vl_logic_vector;
        axi_rd_rresp_c_p4: in     vl_logic_vector(1 downto 0);
        axi_rd_rvalid_c_p4: in     vl_logic;
        axi_rd_data_c_p4: in     vl_logic_vector;
        axi_rd_last_c_p4: in     vl_logic;
        axi_rd_rready_c_p4: out    vl_logic;
        axi_wready_c_p5 : in     vl_logic;
        axi_wid_c_p5    : out    vl_logic_vector;
        axi_waddr_c_p5  : out    vl_logic_vector;
        axi_wlen_c_p5   : out    vl_logic_vector(7 downto 0);
        axi_wsize_c_p5  : out    vl_logic_vector(2 downto 0);
        axi_wburst_c_p5 : out    vl_logic_vector(1 downto 0);
        axi_wlock_c_p5  : out    vl_logic;
        axi_wcache_c_p5 : out    vl_logic_vector(3 downto 0);
        axi_wprot_c_p5  : out    vl_logic_vector(2 downto 0);
        axi_wvalid_c_p5 : out    vl_logic;
        axi_wd_wready_c_p5: in     vl_logic;
        axi_wd_wid_c_p5 : out    vl_logic_vector;
        axi_wd_data_c_p5: out    vl_logic_vector;
        axi_wd_strb_c_p5: out    vl_logic_vector;
        axi_wd_last_c_p5: out    vl_logic;
        axi_wd_valid_c_p5: out    vl_logic;
        axi_wd_bid_c_p5 : in     vl_logic_vector;
        axi_wd_bresp_c_p5: in     vl_logic_vector(1 downto 0);
        axi_wd_bvalid_c_p5: in     vl_logic;
        axi_wd_bready_c_p5: out    vl_logic;
        axi_rready_c_p5 : in     vl_logic;
        axi_rid_c_p5    : out    vl_logic_vector;
        axi_raddr_c_p5  : out    vl_logic_vector;
        axi_rlen_c_p5   : out    vl_logic_vector(7 downto 0);
        axi_rsize_c_p5  : out    vl_logic_vector(2 downto 0);
        axi_rburst_c_p5 : out    vl_logic_vector(1 downto 0);
        axi_rlock_c_p5  : out    vl_logic;
        axi_rcache_c_p5 : out    vl_logic_vector(3 downto 0);
        axi_rprot_c_p5  : out    vl_logic_vector(2 downto 0);
        axi_rvalid_c_p5 : out    vl_logic;
        axi_rd_bid_c_p5 : in     vl_logic_vector;
        axi_rd_rresp_c_p5: in     vl_logic_vector(1 downto 0);
        axi_rd_rvalid_c_p5: in     vl_logic;
        axi_rd_data_c_p5: in     vl_logic_vector;
        axi_rd_last_c_p5: in     vl_logic;
        axi_rd_rready_c_p5: out    vl_logic;
        cmd_err         : out    vl_logic;
        data_msmatch_err: out    vl_logic;
        write_err       : out    vl_logic;
        read_err        : out    vl_logic;
        test_cmptd      : out    vl_logic;
        cmptd_one_wr_rd : out    vl_logic;
        dbg_wr_sts_vld  : out    vl_logic;
        dbg_wr_sts      : out    vl_logic_vector;
        dbg_rd_sts_vld  : out    vl_logic;
        dbg_rd_sts      : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of C_PORT_CONFIG : constant is 1;
    attribute mti_svvh_generic_type of C_P0_PORT_MODE : constant is 1;
    attribute mti_svvh_generic_type of C_P1_PORT_MODE : constant is 1;
    attribute mti_svvh_generic_type of C_P2_PORT_MODE : constant is 1;
    attribute mti_svvh_generic_type of C_P3_PORT_MODE : constant is 1;
    attribute mti_svvh_generic_type of C_P4_PORT_MODE : constant is 1;
    attribute mti_svvh_generic_type of C_P5_PORT_MODE : constant is 1;
    attribute mti_svvh_generic_type of C_PORT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of C_BEGIN_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of C_END_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of C_PRBS_EADDR_MASK_POS : constant is 1;
    attribute mti_svvh_generic_type of C_PRBS_SADDR_MASK_POS : constant is 1;
    attribute mti_svvh_generic_type of C_EN_UPSIZER : constant is 1;
    attribute mti_svvh_generic_type of C_AXI_NBURST_SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of C_ENFORCE_RD_WR : constant is 1;
    attribute mti_svvh_generic_type of C_ENFORCE_RD_WR_CMD : constant is 1;
    attribute mti_svvh_generic_type of C_ENFORCE_RD_WR_PATTERN : constant is 1;
    attribute mti_svvh_generic_type of C_EN_WRAP_TRANS : constant is 1;
    attribute mti_svvh_generic_type of C_P0_AXI_SUPPORTS_READ : constant is 1;
    attribute mti_svvh_generic_type of C_P0_AXI_SUPPORTS_WRITE : constant is 1;
    attribute mti_svvh_generic_type of C_P0_AXI_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P0_AXI_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P0_AXI_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P1_AXI_SUPPORTS_READ : constant is 1;
    attribute mti_svvh_generic_type of C_P1_AXI_SUPPORTS_WRITE : constant is 1;
    attribute mti_svvh_generic_type of C_P1_AXI_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P1_AXI_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P1_AXI_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P2_AXI_SUPPORTS_READ : constant is 1;
    attribute mti_svvh_generic_type of C_P2_AXI_SUPPORTS_WRITE : constant is 1;
    attribute mti_svvh_generic_type of C_P2_AXI_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P2_AXI_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P2_AXI_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P3_AXI_SUPPORTS_READ : constant is 1;
    attribute mti_svvh_generic_type of C_P3_AXI_SUPPORTS_WRITE : constant is 1;
    attribute mti_svvh_generic_type of C_P3_AXI_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P3_AXI_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P3_AXI_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P4_AXI_SUPPORTS_READ : constant is 1;
    attribute mti_svvh_generic_type of C_P4_AXI_SUPPORTS_WRITE : constant is 1;
    attribute mti_svvh_generic_type of C_P4_AXI_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P4_AXI_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P4_AXI_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P5_AXI_SUPPORTS_READ : constant is 1;
    attribute mti_svvh_generic_type of C_P5_AXI_SUPPORTS_WRITE : constant is 1;
    attribute mti_svvh_generic_type of C_P5_AXI_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P5_AXI_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_P5_AXI_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DBG_WR_STS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DBG_RD_STS_WIDTH : constant is 1;
end s6_axi4_tg;
