library verilog;
use verilog.vl_types.all;
entity scrambler_tb is
end scrambler_tb;
